module assign_module (input [3:0] in, output F);
    
endmodule