module counter(input clk, input wire rstn, input [3:0] in, output reg[4:0] out);

