module vector_tb;

reg reset = 0;
reg clk = 0;
wire[3:0]